
-----------------------------------

----- WORD SETUP -----
with binary_select select binary_word(127) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(126) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(125) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(124) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(123) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(122) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(121) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(120) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(119) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(118) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(117) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(116) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(115) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(114) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(113) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(112) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(111) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(110) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(109) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(108) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(107) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(106) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(105) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(104) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(103) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(102) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(101) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(100) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(99) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(98) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(97) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(96) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(95) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(94) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(93) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(92) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(91) <= 
	'0' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(90) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(89) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(88) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(87) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(86) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(85) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(84) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(83) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(82) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(81) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(80) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(79) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(78) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(77) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(76) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(75) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(74) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(73) <= 
	'0' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(72) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(71) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(70) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(69) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(68) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(67) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(66) <= 
	'0' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(65) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(64) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(63) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(62) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(61) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(60) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(59) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(58) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(57) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(56) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(55) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(54) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(53) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(52) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(51) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(50) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(49) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(48) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(47) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(46) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(45) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(44) <= 
	'0' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(43) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(42) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(41) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(40) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(39) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(38) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(37) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(36) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(35) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(34) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(33) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(32) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(31) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(30) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(29) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(28) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(27) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(26) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(25) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(24) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(23) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(22) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(21) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(20) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(19) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(18) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(17) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(16) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(15) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(14) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(13) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(12) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(11) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(10) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(9) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(8) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(7) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(6) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(5) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_word(4) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(3) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(2) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(1) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_word(0) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

-----------------------------------

----- TIP SETUP -----
with binary_select select binary_tip(127) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(126) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(125) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(124) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(123) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(122) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(121) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(120) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(119) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(118) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(117) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(116) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(115) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(114) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(113) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(112) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(111) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(110) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(109) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(108) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(107) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(106) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(105) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(104) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(103) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(102) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(101) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(100) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(99) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(98) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(97) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(96) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(95) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(94) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(93) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(92) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(91) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(90) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(89) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(88) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(87) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(86) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(85) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(84) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(83) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(82) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(81) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(80) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(79) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(78) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(77) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(76) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(75) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(74) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(73) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(72) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(71) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(70) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(69) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(68) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(67) <= 
	'1' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(66) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(65) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(64) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(63) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(62) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(61) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(60) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(59) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(58) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'0' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(57) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(56) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(55) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(54) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(53) <= 
	'0' when "0000000",
	'1' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(52) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(51) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'1' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(50) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'1' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(49) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(48) <= 
	'1' when "0000000",
	'0' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'1' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(47) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(46) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(45) <= 
	'0' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'0' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'1' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'1' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'1' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(44) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(43) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(42) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(41) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(40) <= 
	'1' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'1' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'0' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'0' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'0' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(39) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(38) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(37) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'1' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'0' when "0010101",
	'1' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'0' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'1' when "1000100",
	'0' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'0' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'0' when "1010001",
	'1' when "1010010",
	'0' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'0' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'0' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'0' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'0' when "1101001",
	'1' when "1101010",
	'0' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'0' when "1110001",
	'1' when "1110010",
	'0' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'0' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(36) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(35) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(34) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(33) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'1' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'1' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'1' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(32) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'1' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'1' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'0' when "1000100",
	'1' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'1' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'1' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'1' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'1' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'1' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'1' when "1101001",
	'0' when "1101010",
	'1' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'1' when "1110001",
	'0' when "1110010",
	'1' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'1' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(31) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(30) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(29) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'0' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'0' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'0' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'0' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'0' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'0' when "1111000",
	'1' when "1111001",
	'0' when "1111010",
	'1' when "1111011",
	'0' when "1111100",
	'1' when "1111101",
	'0' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(28) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(27) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(26) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(25) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'1' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'0' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(24) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'1' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'1' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'1' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'1' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'1' when "1111000",
	'0' when "1111001",
	'1' when "1111010",
	'0' when "1111011",
	'1' when "1111100",
	'0' when "1111101",
	'1' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(23) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(22) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(21) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'0' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'0' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'0' when "0101110",
	'1' when "0101111",
	'0' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'0' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(20) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(19) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(18) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(17) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(16) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'1' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'1' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'1' when "0101110",
	'0' when "0101111",
	'1' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'1' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(15) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(14) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(13) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'0' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'0' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(12) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(11) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(10) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(9) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(8) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'1' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'1' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(7) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(6) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(5) <= 
	'1' when "0000000",
	'1' when "0000001",
	'1' when "0000010",
	'1' when "0000011",
	'1' when "0000100",
	'1' when "0000101",
	'1' when "0000110",
	'1' when "0000111",
	'1' when "0001000",
	'1' when "0001001",
	'1' when "0001010",
	'1' when "0001011",
	'1' when "0001100",
	'1' when "0001101",
	'1' when "0001110",
	'1' when "0001111",
	'1' when "0010000",
	'1' when "0010001",
	'1' when "0010010",
	'1' when "0010011",
	'1' when "0010100",
	'1' when "0010101",
	'1' when "0010110",
	'1' when "0010111",
	'1' when "0011000",
	'1' when "0011001",
	'1' when "0011010",
	'1' when "0011011",
	'1' when "0011100",
	'1' when "0011101",
	'1' when "0011110",
	'1' when "0011111",
	'1' when "0100000",
	'1' when "0100001",
	'1' when "0100010",
	'1' when "0100011",
	'1' when "0100100",
	'1' when "0100101",
	'1' when "0100110",
	'1' when "0100111",
	'1' when "0101000",
	'1' when "0101001",
	'1' when "0101010",
	'1' when "0101011",
	'1' when "0101100",
	'1' when "0101101",
	'1' when "0101110",
	'1' when "0101111",
	'1' when "0110000",
	'1' when "0110001",
	'1' when "0110010",
	'1' when "0110011",
	'1' when "0110100",
	'1' when "0110101",
	'1' when "0110110",
	'1' when "0110111",
	'1' when "0111000",
	'1' when "0111001",
	'1' when "0111010",
	'1' when "0111011",
	'1' when "0111100",
	'1' when "0111101",
	'1' when "0111110",
	'1' when "0111111",
	'1' when "1000000",
	'1' when "1000001",
	'1' when "1000010",
	'1' when "1000011",
	'1' when "1000100",
	'1' when "1000101",
	'1' when "1000110",
	'1' when "1000111",
	'1' when "1001000",
	'1' when "1001001",
	'1' when "1001010",
	'1' when "1001011",
	'1' when "1001100",
	'1' when "1001101",
	'1' when "1001110",
	'1' when "1001111",
	'1' when "1010000",
	'1' when "1010001",
	'1' when "1010010",
	'1' when "1010011",
	'1' when "1010100",
	'1' when "1010101",
	'1' when "1010110",
	'1' when "1010111",
	'1' when "1011000",
	'1' when "1011001",
	'1' when "1011010",
	'1' when "1011011",
	'1' when "1011100",
	'1' when "1011101",
	'1' when "1011110",
	'1' when "1011111",
	'1' when "1100000",
	'1' when "1100001",
	'1' when "1100010",
	'1' when "1100011",
	'1' when "1100100",
	'1' when "1100101",
	'1' when "1100110",
	'1' when "1100111",
	'1' when "1101000",
	'1' when "1101001",
	'1' when "1101010",
	'1' when "1101011",
	'1' when "1101100",
	'1' when "1101101",
	'1' when "1101110",
	'1' when "1101111",
	'1' when "1110000",
	'1' when "1110001",
	'1' when "1110010",
	'1' when "1110011",
	'1' when "1110100",
	'1' when "1110101",
	'1' when "1110110",
	'1' when "1110111",
	'1' when "1111000",
	'1' when "1111001",
	'1' when "1111010",
	'1' when "1111011",
	'1' when "1111100",
	'1' when "1111101",
	'1' when "1111110",
	'1' when "1111111",
	'0' when others;

with binary_select select binary_tip(4) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(3) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(2) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(1) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

with binary_select select binary_tip(0) <= 
	'0' when "0000000",
	'0' when "0000001",
	'0' when "0000010",
	'0' when "0000011",
	'0' when "0000100",
	'0' when "0000101",
	'0' when "0000110",
	'0' when "0000111",
	'0' when "0001000",
	'0' when "0001001",
	'0' when "0001010",
	'0' when "0001011",
	'0' when "0001100",
	'0' when "0001101",
	'0' when "0001110",
	'0' when "0001111",
	'0' when "0010000",
	'0' when "0010001",
	'0' when "0010010",
	'0' when "0010011",
	'0' when "0010100",
	'0' when "0010101",
	'0' when "0010110",
	'0' when "0010111",
	'0' when "0011000",
	'0' when "0011001",
	'0' when "0011010",
	'0' when "0011011",
	'0' when "0011100",
	'0' when "0011101",
	'0' when "0011110",
	'0' when "0011111",
	'0' when "0100000",
	'0' when "0100001",
	'0' when "0100010",
	'0' when "0100011",
	'0' when "0100100",
	'0' when "0100101",
	'0' when "0100110",
	'0' when "0100111",
	'0' when "0101000",
	'0' when "0101001",
	'0' when "0101010",
	'0' when "0101011",
	'0' when "0101100",
	'0' when "0101101",
	'0' when "0101110",
	'0' when "0101111",
	'0' when "0110000",
	'0' when "0110001",
	'0' when "0110010",
	'0' when "0110011",
	'0' when "0110100",
	'0' when "0110101",
	'0' when "0110110",
	'0' when "0110111",
	'0' when "0111000",
	'0' when "0111001",
	'0' when "0111010",
	'0' when "0111011",
	'0' when "0111100",
	'0' when "0111101",
	'0' when "0111110",
	'0' when "0111111",
	'0' when "1000000",
	'0' when "1000001",
	'0' when "1000010",
	'0' when "1000011",
	'0' when "1000100",
	'0' when "1000101",
	'0' when "1000110",
	'0' when "1000111",
	'0' when "1001000",
	'0' when "1001001",
	'0' when "1001010",
	'0' when "1001011",
	'0' when "1001100",
	'0' when "1001101",
	'0' when "1001110",
	'0' when "1001111",
	'0' when "1010000",
	'0' when "1010001",
	'0' when "1010010",
	'0' when "1010011",
	'0' when "1010100",
	'0' when "1010101",
	'0' when "1010110",
	'0' when "1010111",
	'0' when "1011000",
	'0' when "1011001",
	'0' when "1011010",
	'0' when "1011011",
	'0' when "1011100",
	'0' when "1011101",
	'0' when "1011110",
	'0' when "1011111",
	'0' when "1100000",
	'0' when "1100001",
	'0' when "1100010",
	'0' when "1100011",
	'0' when "1100100",
	'0' when "1100101",
	'0' when "1100110",
	'0' when "1100111",
	'0' when "1101000",
	'0' when "1101001",
	'0' when "1101010",
	'0' when "1101011",
	'0' when "1101100",
	'0' when "1101101",
	'0' when "1101110",
	'0' when "1101111",
	'0' when "1110000",
	'0' when "1110001",
	'0' when "1110010",
	'0' when "1110011",
	'0' when "1110100",
	'0' when "1110101",
	'0' when "1110110",
	'0' when "1110111",
	'0' when "1111000",
	'0' when "1111001",
	'0' when "1111010",
	'0' when "1111011",
	'0' when "1111100",
	'0' when "1111101",
	'0' when "1111110",
	'0' when "1111111",
	'0' when others;

-----------------------------------
