library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity banco_lvl3 is
	port(
        binary_select: in std_logic_vector(5 downto 0);
        binary_tip : out std_logic_vector(127 downto 0);
        binary_word : out std_logic_vector(127 downto 0)
    );
end entity;

architecture arch_banco_lvl3 of banco_lvl3 is
    begin

-----------------------------------

----- WORD SETUP -----
with binary_select select binary_word(127) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(126) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(125) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(124) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(123) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(122) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(121) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(120) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(119) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(118) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(117) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(116) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(115) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(114) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(113) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(112) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(111) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(110) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(109) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(108) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(107) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(106) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(105) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(104) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(103) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(102) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(101) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(100) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(99) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(98) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(97) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(96) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(95) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(94) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(93) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(92) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(91) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(90) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(89) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(88) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(87) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(86) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(85) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(84) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(83) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(82) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(81) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(80) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(79) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(78) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(77) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(76) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(75) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(74) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(73) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(72) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(71) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(70) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(69) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(68) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(67) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(66) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(65) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(64) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(63) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(62) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(61) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(60) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(59) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(58) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(57) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(56) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(55) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(54) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(53) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(52) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(51) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(50) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(49) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(48) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(47) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(46) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(45) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(44) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(43) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(42) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(41) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(40) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(39) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(38) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(37) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(36) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(35) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(34) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(33) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(32) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(31) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(30) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(29) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(28) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(27) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(26) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(25) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(24) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(23) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(22) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(21) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(20) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(19) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(18) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(17) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(16) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(15) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(14) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(13) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(12) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(11) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(10) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(9) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(8) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(7) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(6) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(5) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(4) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_word(3) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(2) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(1) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_word(0) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

-----------------------------------

----- TIP SETUP -----
with binary_select select binary_tip(127) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(126) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(125) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(124) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(123) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(122) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(121) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(120) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(119) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(118) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(117) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(116) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(115) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(114) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(113) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(112) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(111) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(110) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(109) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(108) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(107) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(106) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(105) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(104) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(103) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(102) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(101) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(100) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(99) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(98) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(97) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(96) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(95) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(94) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(93) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(92) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(91) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(90) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(89) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(88) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(87) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(86) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(85) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(84) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(83) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(82) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(81) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(80) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(79) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(78) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(77) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(76) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(75) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(74) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(73) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(72) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(71) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(70) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(69) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(68) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(67) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(66) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(65) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(64) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(63) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(62) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(61) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(60) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(59) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(58) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(57) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(56) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(55) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(54) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(53) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(52) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(51) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(50) <=
	'1' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(49) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(48) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(47) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(46) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(45) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(44) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(43) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(42) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(41) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(40) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(39) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(38) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(37) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(36) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(35) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(34) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'1' when "100100",
	'0' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(33) <=
	'0' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(32) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'1' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'1' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(31) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(30) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(29) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(28) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'1' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(27) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(26) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'1' when "001011",
	'0' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(25) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'0' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'1' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(24) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'0' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'0' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(23) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(22) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(21) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(20) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'0' when "010111",
	'0' when "011000",
	'1' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(19) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'0' when "000011",
	'0' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'1' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(18) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(17) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'1' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(16) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'0' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(15) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(14) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(13) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(12) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'0' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(11) <=
	'0' when "000000",
	'1' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'1' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'0' when "011001",
	'1' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'1' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'1' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'1' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'1' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(10) <=
	'1' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'1' when "001011",
	'0' when "001100",
	'0' when "001101",
	'1' when "001110",
	'0' when "001111",
	'1' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'1' when "011101",
	'1' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'0' when "100110",
	'1' when "100111",
	'0' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'0' when "111000",
	'1' when "111001",
	'0' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(9) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'1' when "110010",
	'0' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(8) <=
	'0' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'0' when "001011",
	'1' when "001100",
	'1' when "001101",
	'0' when "001110",
	'1' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'1' when "010011",
	'0' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'0' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'1' when "100110",
	'0' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'0' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'1' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(7) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(6) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'1' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(5) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'0' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'0' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(4) <=
	'0' when "000000",
	'0' when "000001",
	'0' when "000010",
	'0' when "000011",
	'0' when "000100",
	'0' when "000101",
	'0' when "000110",
	'0' when "000111",
	'0' when "001000",
	'0' when "001001",
	'0' when "001010",
	'0' when "001011",
	'0' when "001100",
	'0' when "001101",
	'0' when "001110",
	'0' when "001111",
	'0' when "010000",
	'1' when "010001",
	'0' when "010010",
	'0' when "010011",
	'0' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'0' when "011000",
	'0' when "011001",
	'0' when "011010",
	'0' when "011011",
	'0' when "011100",
	'0' when "011101",
	'0' when "011110",
	'0' when "011111",
	'1' when "100000",
	'0' when "100001",
	'0' when "100010",
	'0' when "100011",
	'0' when "100100",
	'0' when "100101",
	'0' when "100110",
	'0' when "100111",
	'0' when "101000",
	'0' when "101001",
	'0' when "101010",
	'0' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'0' when "110000",
	'0' when "110001",
	'0' when "110010",
	'0' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'0' when "110111",
	'0' when "111000",
	'0' when "111001",
	'0' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'0' when "111110",
	'0' when "111111",
	'0' when others;

with binary_select select binary_tip(3) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'0' when "101101",
	'1' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(2) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'1' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'0' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'1' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'0' when "100000",
	'1' when "100001",
	'0' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'0' when "101010",
	'1' when "101011",
	'1' when "101100",
	'1' when "101101",
	'1' when "101110",
	'1' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'1' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(1) <=
	'1' when "000000",
	'0' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'0' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'0' when "010011",
	'1' when "010100",
	'0' when "010101",
	'0' when "010110",
	'0' when "010111",
	'1' when "011000",
	'1' when "011001",
	'0' when "011010",
	'1' when "011011",
	'1' when "011100",
	'0' when "011101",
	'0' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'0' when "100010",
	'0' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'0' when "101001",
	'0' when "101010",
	'1' when "101011",
	'0' when "101100",
	'0' when "101101",
	'0' when "101110",
	'0' when "101111",
	'1' when "110000",
	'0' when "110001",
	'1' when "110010",
	'1' when "110011",
	'0' when "110100",
	'0' when "110101",
	'0' when "110110",
	'1' when "110111",
	'1' when "111000",
	'0' when "111001",
	'1' when "111010",
	'0' when "111011",
	'0' when "111100",
	'1' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;

with binary_select select binary_tip(0) <=
	'1' when "000000",
	'1' when "000001",
	'1' when "000010",
	'1' when "000011",
	'1' when "000100",
	'0' when "000101",
	'1' when "000110",
	'1' when "000111",
	'1' when "001000",
	'1' when "001001",
	'1' when "001010",
	'1' when "001011",
	'1' when "001100",
	'1' when "001101",
	'1' when "001110",
	'1' when "001111",
	'1' when "010000",
	'1' when "010001",
	'1' when "010010",
	'1' when "010011",
	'1' when "010100",
	'0' when "010101",
	'1' when "010110",
	'1' when "010111",
	'1' when "011000",
	'1' when "011001",
	'1' when "011010",
	'1' when "011011",
	'1' when "011100",
	'1' when "011101",
	'1' when "011110",
	'1' when "011111",
	'1' when "100000",
	'1' when "100001",
	'1' when "100010",
	'1' when "100011",
	'1' when "100100",
	'1' when "100101",
	'1' when "100110",
	'1' when "100111",
	'1' when "101000",
	'1' when "101001",
	'1' when "101010",
	'1' when "101011",
	'0' when "101100",
	'1' when "101101",
	'0' when "101110",
	'1' when "101111",
	'1' when "110000",
	'1' when "110001",
	'1' when "110010",
	'1' when "110011",
	'1' when "110100",
	'0' when "110101",
	'1' when "110110",
	'1' when "110111",
	'1' when "111000",
	'1' when "111001",
	'1' when "111010",
	'1' when "111011",
	'1' when "111100",
	'0' when "111101",
	'1' when "111110",
	'1' when "111111",
	'0' when others;
-----------------------------------
end architecture;