library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity word_selector is
    port(
        data_in : in std_logic_vector(1 downto 0);
        data_out : out std_logic_vector(255 downto 0)
    );
end entity;

architecture behav of word_selector is
    begin
        data_out <=
            "0000100000100000001000000101001001000101010001110100100101010011" &
            "0101010001010010010000010100010001001111010100100010000000100000" &
            "0010000000100000001000000100001101101111011011010111000001101111" &
            "0110111001100101011011100111010001100101001000000010000000100000" when data_in = "01" else

            "0010000000100000001000000100101001010101010000100100100101001100" &
            "0100000101001101010001010100111001010100010011110010000000100000" &
            "0010000000100000001000000010000000100000010100000111010101101110" &
            "0110100101100011011000010110111100100000001000000010000000100000" when data_in = "10" else

            "0100011001000101010011000100100101010000010001010010000001010110" &
            "0100000101001100010001010100111001000011010010010100000100100000" &
            "0010000000100000010100010111010101100101001000000110001101100001" &
            "0111001001100001001000000110001001101111011011010010000000100000" when data_in = "11" else
            
            "0000000000000000000000000000000000000000000000000000000000000000" &
            "0000000000000000000000000000000000000000000000000000000000000000" &
            "0000000000000000000000000000000000000000000000000000000000000000" &
            "0000000000000000000000000000000000000000000000000000000000000000"; --00

            --00: fácil -> REGISTRADOR / dica: Componente
            --01: médio -> JUBILAMENTO / dica: Punicao
            --11: politécnico -> FELIPE VALENCIA / dica: Que cara bom

end architecture;


