--screens_register1: armazena os códigos ASCII das telas de introdução e dificuldade
library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity screens_register1 is
    port(
        screen_number : in std_logic_vector(1 downto 0);
        code_out : out std_logic_vector(255 downto 0)
    );
end entity;

architecture behav of screens_register1 is
    begin
        code_out <=
            "0010000000100000010010100100111101000111010011110010000001000100" &
            "0100000100100000010001100100111101010010010000110100000100100000" &
            "0010000001100011011010000110010101101001011100100110000100100000" &
            "0110000100100000011100110111010101100011011011110011111100100000" when screen_number = "00" else

            "0010000000100000010001000110100101100110011010010110001101110101" &
            "0110110001100100011000010110010001100101001110100010000000100000" &
            "0011110000101101001000000010000000100000001000000100011001100001" &
            "0110001101101001011011000010000000100000001000000010110100111110" when screen_number = "01" else

            "0010000000100000010001000110100101100110011010010110001101110101" &
            "0110110001100100011000010110010001100101001110100010000000100000" &
            "0011110000101101001000000010000000100000001000000100110101100101" &
            "0110010001101001011011110010000000100000001000000010110100111110" when screen_number = "10" else

            "0010000000100000010001000110100101100110011010010110001101110101" &
            "0110110001100100011000010110010001100101001110100010000000100000" &
            "0011110000101101001000000101000001101111011011000110100101110100" &
            "0110010101100011011011100110100101100011011011110010110100111110"; --when screen_number = "11"


            -- "00" :
            -- JOGO DA FORCA
            -- cheira a suco?

            -- "01" : 
            -- Dificuldade:
            -- <- Facil ->

            --  "10" : 
            -- Dificuldade:
            -- <- Medio ->

            -- "11" :
            -- Dificuldade:
            -- <-Politecnico->
    end architecture;